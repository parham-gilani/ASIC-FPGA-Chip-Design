library verilog;
use verilog.vl_types.all;
entity Part1_vlg_vec_tst is
end Part1_vlg_vec_tst;
