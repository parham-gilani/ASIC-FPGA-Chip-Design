module handshake_p1(input clock, reset,
					input [3:0] ps2_data, input ts,
					output reg [3:0] leds);

// Your code goes here...

endmodule
