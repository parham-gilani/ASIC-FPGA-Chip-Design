library verilog;
use verilog.vl_types.all;
entity Part3_vlg_vec_tst is
end Part3_vlg_vec_tst;
